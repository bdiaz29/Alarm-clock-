

module project( SW, CLK,  LED,SSEG_AN,SSEG_CA, PBR, PBL);
 output reg [7:0] SSEG_CA;
 output reg [7:0] SSEG_AN;
 //output reg Alarm;
 //input  PBL;
 input  PBR;
 input  PBL;
 //input  PBB;
input[1:0] SW;
input CLK;
output reg [1:0] LED;
reg [2:0] counter;
reg [6:0] second;
reg [6:0] minute;
reg [5:0] hour;

reg [6:0] set_second;
reg [6:0] set_minute;
reg [5:0] set_hour;


reg set_minC;
reg set_HC;
reg min_C;
reg H_C;


always
begin
set_second=0;
//LED[1]=PBL;
end






reg scape;

reg [7:0] temp;
always 
begin
temp=8'd55;
end

reg speed;

always
begin
if((set_hour==hour)&&(set_minute==minute))
begin
LED[0]=1;
end
else
begin
LED[0]=0;
end

end

//display clock
pwmclock P(CLK, pwm_clk);
//refrence clocks
secClk S(CLK,SW[0],secCLK);
minClk M(secCLK,minCLK);
hClk H(min_C,hCLK);
initial
begin
second=0;
minute=0;
hour=0;
set_second=0;
set_minute=0;
set_hour=0;
end

always
begin
case(SW)
1'b0 : 
begin
speed=1'b0;
end
1'b1 :
begin
speed=1'b1;
end

endcase
end
////////////////////////////////////////////////////////
always @(posedge pwm_clk)
begin
counter=counter+1; 
end
//seconds
always @(posedge secCLK)
begin
second=second+1;

case(second)
6'd60 :second=0;
6'd61 :second=0;
6'd62 :second=0;
6'd63 :second=0;
default:second=second;
endcase

end
//hours
always @(posedge H_C)
begin
hour=hour+1;
case(hour)
5'd24:hour=0;
5'd25:hour=0;
5'd26:hour=0;
5'd27:hour=0;
5'd28:hour=0;
5'd29:hour=0;
5'd30:hour=0;
default:hour=hour;
endcase
end

always
begin
H_C=hCLK|(PBL&(~SW[1]));
//H_C=0;
set_HC=PBL&SW[1];
end

always@(posedge set_HC)
begin
set_hour=set_hour+1;
case(set_hour)
5'd24:set_hour=0;
5'd25:set_hour=0;
5'd26:set_hour=0;
5'd27:set_hour=0;
5'd28:set_hour=0;
5'd29:set_hour=0;
5'd30:set_hour=0;
default:set_hour=set_hour;
endcase
end



always @(posedge min_C)
begin
minute=minute+1;
case(minute)
6'd60:minute=0;
6'd61:minute=0;
6'd62:minute=0;
6'd63:minute=0;
default:minute=minute;
endcase


end

always@(posedge set_minC)
begin
set_minute=set_minute+1;
case(set_minute)
6'd59:set_minute=0;
6'd60:set_minute=0;
6'd61:set_minute=0;
6'd62:set_minute=0;
6'd63:set_minute=0;
default:set_minute=set_minute;
endcase
end

always
begin
min_C=minCLK|(PBR&(~SW[1]));
set_minC=PBR&SW[1];
end
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////



always 
begin
case(SW[1])
1'b0:
begin
///////////////////////////////////////////////
case(counter)
//lower second
3'd0:begin
case(second)//lower bound second
6'd0:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd1:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd2:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd3:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd4:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd5:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd6:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd7:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd8:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd9:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd10:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd11:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd13:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd14:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd15:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd16:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd17:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd18:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd19:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd20:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd21:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd22:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd24:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd25:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd26:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd27:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd28:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd29:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd30:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd31:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd32:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd33:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd34:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd35:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd36:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd37:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd38:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd39:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd40:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd41:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd42:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd43:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd44:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd45:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd46:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd47:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd48:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd49:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd50:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd51:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd52:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd53:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd54:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd55:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd56:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd57:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd58:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd59:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd60:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
default:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
endcase
end
3'd1:begin
case(second)//upper bound second
6'd0:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end//0
6'd1:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///1
6'd2:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///2
6'd3:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///3
6'd4:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///4
6'd5:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///5
6'd6:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///6
6'd7:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///7
6'd8:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///8
6'd9:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///9
6'd10:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end//1
6'd11:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd13:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd14:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd15:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd16:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd17:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd18:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd19:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd20:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end//2
6'd21:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd22:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd24:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd25:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd26:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd27:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd28:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd29:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd30:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end//3
6'd31:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd32:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd33:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd34:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd35:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd36:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd37:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd38:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd39:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd40:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end//4
6'd41:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd42:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd43:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd44:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd45:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd46:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd47:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd48:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd49:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd50:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end//5
6'd51:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd52:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd53:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd54:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd55:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd56:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd57:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd58:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd59:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd60:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10000010;end//6
default:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end//0
endcase
end
3'd2:begin
case(minute)//minute lower bound
6'd0:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd1:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd2:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd3:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd4:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd5:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd6:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd7:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd8:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd9:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd10:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd11:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd13:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd14:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd15:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd16:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd17:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd18:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd19:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd20:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd21:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd22:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd24:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd25:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd26:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd27:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd28:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd29:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd30:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd31:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd32:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd33:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd34:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd35:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd36:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd37:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd38:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd39:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd40:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd41:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd42:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd43:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd44:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd45:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd46:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd47:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd48:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd49:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd50:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd51:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd52:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd53:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd54:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd55:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd56:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd57:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd58:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd59:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd60:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
default:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
endcase
end
3'd3:begin
case(minute)//minute upper bound
6'd0:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end//0
6'd1:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///1
6'd2:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///2
6'd3:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///3
6'd4:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///4
6'd5:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///5
6'd6:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///6
6'd7:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///7
6'd8:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///8
6'd9:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///9
6'd10:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end//1
6'd11:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd13:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd14:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd15:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd16:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd17:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd18:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd19:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd20:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end//2
6'd21:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd22:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd24:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd25:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd26:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd27:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd28:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd29:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd30:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end//3
6'd31:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd32:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd33:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd34:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd35:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd36:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd37:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd38:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd39:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd40:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end//4
6'd41:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd42:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd43:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd44:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd45:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd46:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd47:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd48:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd49:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd50:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end//5
6'd51:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd52:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd53:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd54:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd55:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd56:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd57:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd58:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd59:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd60:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10000010;end//6
default:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end//0
endcase
end
3'd4:begin
case(hour)//hour lower bound
6'd0:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11000000;end
6'd1:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11111001;end
6'd2:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10100100;end
6'd3:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10110000;end
6'd4:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10011001;end
6'd5:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10010010;end
6'd6:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10000010;end
6'd7:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11111000;end
6'd8:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10000000;end
6'd9:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10010000;end
6'd10:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11000000;end
6'd11:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10100100;end
6'd13:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10110000;end
6'd14:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10011001;end
6'd15:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10010010;end
6'd16:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10000010;end
6'd17:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11111000;end
6'd18:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10000000;end
6'd19:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10010000;end
6'd20:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11000000;end
6'd21:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11111001;end
6'd22:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10110000;end
6'd24:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10011001;end
default:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11000000;end
endcase
end
3'd5:begin
case(hour)//set hour upper bound
6'd0:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end//0
6'd1:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///1
6'd2:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///2
6'd3:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///3
6'd4:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///4
6'd5:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///5
6'd6:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///6
6'd7:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///7
6'd8:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///8
6'd9:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///9
6'd10:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end//1
6'd11:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd13:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd14:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd15:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd16:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd17:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd18:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd19:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd20:begin SSEG_AN=8'b11011111;SSEG_CA=8'b10100100;end//2
6'd21:begin SSEG_AN=8'b11011111;SSEG_CA=8'b10100100;end
6'd22:begin SSEG_AN=8'b11011111;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11011111;SSEG_CA=8'b10100100;end
6'd24:begin SSEG_AN=8'b11011111;SSEG_CA=8'b10100100;end
default:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end//0
endcase
end
3'd6:
begin
case(temp)//temp lower bound
8'd0:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd1:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd2:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd3:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd4:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd5:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd6:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd7:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd8:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd9:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd10:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd11:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd12:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd13:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd14:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd15:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd16:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd17:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd18:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd19:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd20:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd21:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd22:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd23:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd24:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd25:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd26:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd27:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd28:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd29:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd30:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd31:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd32:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd33:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd34:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd35:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd36:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd37:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd38:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd39:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd40:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd41:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd42:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd43:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd44:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd45:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd46:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd47:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd48:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd49:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd50:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd51:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd52:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd53:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd54:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd55:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd56:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd57:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd58:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd59:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd60:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd61:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd62:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd63:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd64:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd65:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd66:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd67:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd68:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd69:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd70:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd71:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd72:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd73:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd74:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd75:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd76:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd77:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd78:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd79:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd80:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd81:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd82:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd83:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd84:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd85:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd86:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd87:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd88:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd89:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd90:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd91:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd92:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd93:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd94:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd95:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd96:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd97:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd98:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd99:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
default:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
endcase
end
//temp upper bound
3'd7:
begin
case(temp)//temp upper bound
8'd0:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end//0
8'd1:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///1
8'd2:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///2
8'd3:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///3
8'd4:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///4
8'd5:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///5
8'd6:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///6
8'd7:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///7
8'd8:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///8
8'd9:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///9
8'd10:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end//1
8'd11:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd12:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd13:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd14:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd15:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd16:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd17:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd18:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd19:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd20:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end//2
8'd21:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd22:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd23:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd24:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd25:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd26:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd27:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd28:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd29:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd30:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end//3
8'd31:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd32:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd33:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd34:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd35:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd36:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd37:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd38:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd39:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd40:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end//4
8'd41:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd42:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd43:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd44:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd45:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd46:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd47:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd48:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd49:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd50:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end//5
8'd51:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd52:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd53:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd54:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd55:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd56:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd57:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd58:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd59:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd60:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end//6
8'd61:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end//0
8'd62:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd63:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd64:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd65:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd66:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd67:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd68:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd69:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd70:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end//7
8'd71:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd72:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd73:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd74:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd75:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd76:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd77:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd78:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd79:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd80:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end///8
8'd81:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd82:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd83:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd84:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd85:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd86:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd87:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd88:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd89:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd90:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end//9
8'd91:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd92:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd93:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd94:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd95:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd96:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd97:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd98:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd99:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
default:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end//0
endcase
end
endcase
///////////////////////////////////////////////
end
1'b1:
begin
//////////////////////////////////////////////
case(counter)
//lower second
3'd0:begin
case(set_second)//lower bound second
6'd0:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd1:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd2:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd3:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd4:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd5:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd6:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd7:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd8:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd9:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd10:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd11:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd13:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd14:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd15:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd16:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd17:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd18:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd19:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd20:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd21:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd22:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd24:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd25:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd26:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd27:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd28:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd29:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd30:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd31:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd32:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd33:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd34:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd35:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd36:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd37:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd38:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd39:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd40:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd41:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd42:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd43:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd44:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd45:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd46:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd47:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd48:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd49:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd50:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
6'd51:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111001;end
6'd52:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10100100;end
6'd53:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10110000;end
6'd54:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10011001;end
6'd55:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010010;end
6'd56:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000010;end
6'd57:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11111000;end
6'd58:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10000000;end
6'd59:begin SSEG_AN=8'b11111110;SSEG_CA=8'b10010000;end
6'd60:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
default:begin SSEG_AN=8'b11111110;SSEG_CA=8'b11000000;end
endcase
end
3'd1:begin
case(set_second)//upper bound second
6'd0:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end//0
6'd1:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///1
6'd2:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///2
6'd3:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///3
6'd4:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///4
6'd5:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///5
6'd6:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///6
6'd7:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///7
6'd8:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///8
6'd9:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end///9
6'd10:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end//1
6'd11:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd13:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd14:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd15:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd16:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd17:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd18:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd19:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11111001;end
6'd20:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end//2
6'd21:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd22:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd24:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd25:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd26:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd27:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd28:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd29:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10100100;end
6'd30:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end//3
6'd31:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd32:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd33:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd34:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd35:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd36:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd37:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd38:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd39:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10110000;end
6'd40:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end//4
6'd41:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd42:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd43:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd44:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd45:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd46:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd47:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd48:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd49:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10011001;end
6'd50:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end//5
6'd51:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd52:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd53:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd54:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd55:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd56:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd57:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd58:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd59:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10010010;end
6'd60:begin SSEG_AN=8'b11111101;SSEG_CA=8'b10000010;end//6
default:begin SSEG_AN=8'b11111101;SSEG_CA=8'b11000000;end//0
endcase
end
3'd2:begin
case(set_minute)//minute lower bound
6'd0:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd1:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd2:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd3:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd4:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd5:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd6:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd7:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd8:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd9:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd10:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd11:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd13:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd14:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd15:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd16:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd17:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd18:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd19:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd20:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd21:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd22:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd24:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd25:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd26:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd27:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd28:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd29:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd30:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd31:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd32:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd33:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd34:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd35:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd36:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd37:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd38:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd39:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd40:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd41:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd42:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd43:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd44:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd45:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd46:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd47:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd48:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd49:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd50:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
6'd51:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111001;end
6'd52:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10100100;end
6'd53:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10110000;end
6'd54:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10011001;end
6'd55:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010010;end
6'd56:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000010;end
6'd57:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11111000;end
6'd58:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10000000;end
6'd59:begin SSEG_AN=8'b11111011;SSEG_CA=8'b10010000;end
6'd60:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
default:begin SSEG_AN=8'b11111011;SSEG_CA=8'b11000000;end
endcase
end
3'd3:begin
case(set_minute)//minute upper bound
6'd0:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end//0
6'd1:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///1
6'd2:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///2
6'd3:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///3
6'd4:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///4
6'd5:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///5
6'd6:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///6
6'd7:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///7
6'd8:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///8
6'd9:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end///9
6'd10:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end//1
6'd11:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd13:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd14:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd15:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd16:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd17:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd18:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd19:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11111001;end
6'd20:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end//2
6'd21:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd22:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd24:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd25:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd26:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd27:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd28:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd29:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10100100;end
6'd30:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end//3
6'd31:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd32:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd33:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd34:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd35:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd36:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd37:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd38:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd39:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10110000;end
6'd40:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end//4
6'd41:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd42:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd43:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd44:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd45:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd46:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd47:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd48:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd49:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10011001;end
6'd50:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end//5
6'd51:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd52:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd53:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd54:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd55:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd56:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd57:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd58:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd59:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10010010;end
6'd60:begin SSEG_AN=8'b11110111;SSEG_CA=8'b10000010;end//6
default:begin SSEG_AN=8'b11110111;SSEG_CA=8'b11000000;end//0
endcase
end
3'd4:begin
case(set_hour)//hour lower bound
6'd0:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11000000;end
6'd1:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11111001;end
6'd2:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10100100;end
6'd3:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10110000;end
6'd4:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10011001;end
6'd5:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10010010;end
6'd6:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10000010;end
6'd7:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11111000;end
6'd8:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10000000;end
6'd9:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10010000;end
6'd10:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11000000;end
6'd11:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10100100;end
6'd13:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10110000;end
6'd14:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10011001;end
6'd15:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10010010;end
6'd16:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10000010;end
6'd17:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11111000;end
6'd18:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10000000;end
6'd19:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10010000;end
6'd20:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11000000;end
6'd21:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11111001;end
6'd22:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10110000;end
6'd24:begin SSEG_AN=8'b11101111;SSEG_CA=8'b10011001;end
default:begin SSEG_AN=8'b11101111;SSEG_CA=8'b11000000;end
endcase
end
3'd5:begin
case(set_hour)//set hour upper bound
6'd0:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end//0
6'd1:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///1
6'd2:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///2
6'd3:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///3
6'd4:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///4
6'd5:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///5
6'd6:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///6
6'd7:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///7
6'd8:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///8
6'd9:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end///9
6'd10:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end//1
6'd11:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd12:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd13:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd14:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd15:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd16:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd17:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd18:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd19:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11111001;end
6'd20:begin SSEG_AN=8'b11011111;SSEG_CA=8'b10100100;end//2
6'd21:begin SSEG_AN=8'b11011111;SSEG_CA=8'b10100100;end
6'd22:begin SSEG_AN=8'b11011111;SSEG_CA=8'b10100100;end
6'd23:begin SSEG_AN=8'b11011111;SSEG_CA=8'b10100100;end
6'd24:begin SSEG_AN=8'b11011111;SSEG_CA=8'b10100100;end
default:begin SSEG_AN=8'b11011111;SSEG_CA=8'b11000000;end//0
endcase
end
3'd6:
begin
case(temp)//temp lower bound
8'd0:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd1:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd2:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd3:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd4:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd5:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd6:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd7:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd8:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd9:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd10:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd11:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd12:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd13:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd14:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd15:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd16:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd17:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd18:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd19:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd20:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd21:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd22:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd23:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd24:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd25:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd26:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd27:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd28:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd29:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd30:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd31:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd32:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd33:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd34:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd35:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd36:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd37:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd38:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd39:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd40:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd41:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd42:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd43:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd44:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd45:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd46:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd47:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd48:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd49:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd50:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd51:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd52:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd53:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd54:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd55:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd56:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd57:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd58:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd59:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd60:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd61:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd62:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd63:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd64:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd65:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd66:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd67:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd68:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd69:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd70:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd71:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd72:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd73:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd74:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd75:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd76:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd77:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd78:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd79:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd80:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd81:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd82:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd83:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd84:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd85:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd86:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd87:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd88:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd89:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
8'd90:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010000;end
8'd91:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
8'd92:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111001;end
8'd93:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10100100;end
8'd94:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10110000;end
8'd95:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10011001;end
8'd96:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10010010;end
8'd97:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000010;end
8'd98:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11111000;end
8'd99:begin SSEG_AN=8'b10111111;SSEG_CA=8'b10000000;end
default:begin SSEG_AN=8'b10111111;SSEG_CA=8'b11000000;end
endcase
end
//temp upper bound
3'd7:
begin
case(temp)//temp upper bound
8'd0:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end//0
8'd1:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///1
8'd2:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///2
8'd3:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///3
8'd4:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///4
8'd5:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///5
8'd6:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///6
8'd7:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///7
8'd8:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///8
8'd9:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end///9
8'd10:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end//1
8'd11:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd12:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd13:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd14:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd15:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd16:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd17:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd18:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd19:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111001;end
8'd20:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end//2
8'd21:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd22:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd23:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd24:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd25:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd26:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd27:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd28:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd29:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10100100;end
8'd30:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end//3
8'd31:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd32:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd33:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd34:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd35:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd36:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd37:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd38:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd39:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10110000;end
8'd40:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end//4
8'd41:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd42:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd43:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd44:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd45:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd46:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd47:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd48:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd49:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10011001;end
8'd50:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end//5
8'd51:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd52:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd53:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd54:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd55:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd56:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd57:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd58:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd59:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010010;end
8'd60:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end//6
8'd61:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end//0
8'd62:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd63:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd64:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd65:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd66:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd67:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd68:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd69:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000010;end
8'd70:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end//7
8'd71:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd72:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd73:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd74:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd75:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd76:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd77:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd78:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd79:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11111000;end
8'd80:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end///8
8'd81:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd82:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd83:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd84:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd85:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd86:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd87:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd88:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd89:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10000000;end
8'd90:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end//9
8'd91:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd92:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd93:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd94:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd95:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd96:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd97:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd98:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
8'd99:begin SSEG_AN=8'b01111111;SSEG_CA=8'b10010000;end
default:begin SSEG_AN=8'b01111111;SSEG_CA=8'b11000000;end//0
endcase
end
endcase
//////////////////////////////////////////////
end
endcase
end
//////////////////////////////////////////////////////////////////////
endmodule

//the second clock
//s determines if its running fast or norma;
module secClk(clk,S,secCLK);
input clk;
input S;
reg [31:0] compare;
output reg secCLK;
reg [31:0] counter_out;
	initial begin
	counter_out<= 32'h00000000;
	secCLK <=0;
	end	
	always
	begin
	case(S)
	1'b0:compare=32'h02FAF07F;
	//1'b1:compare=32'h000CB734;
	1'b1:compare=32'h00014585;
	endcase
	end
//this always block runs on the fast 100MHz clock
always @(posedge clk) begin
	counter_out<=    counter_out + 32'h00000001;		
	if (counter_out  > compare) begin 
		counter_out<= 32'h00000000;
		secCLK <= !secCLK;
		end
	end
	
endmodule



///the minute clock
module minClk(clk,minCLK);
input clk;
reg [35:0] counter_out;
reg [35:0] compare;
output reg minCLK;
	initial begin
	counter_out<= 36'h000000000;
	compare=36'h00000003A;
	minCLK <=0;
	end	
//this always block runs on the fast 100MHz clock
always @(posedge clk) begin
	counter_out<=    counter_out + 36'h000000001;		
	if (counter_out  > compare) begin 
		counter_out<= 36'h000000000;
		minCLK <= !minCLK;
		compare=36'h00000001C;
		end
	end

endmodule

///the hour 
module hClk(clk,hCLK);
input clk;
reg [39:0] counter_out;
reg [39:0] compare;
output reg hCLK;
	initial begin
	counter_out<= 40'h0000000000;
	compare=36'h00000003A;
	hCLK <=0;
	end	
//this always block runs on the fast 100MHz clock
always @(posedge clk) begin
	counter_out<=    counter_out + 40'h0000000001;		
	if (counter_out  > compare) begin 
		counter_out<= 40'h0000000000;
		hCLK <= !hCLK;
		compare=40'h000000001C;
		end
	end

endmodule

//500 hz clock
module pwmclock(clk, pwm_clk);
input clk;
reg [31:0] counter_out;
output reg pwm_clk;
	initial begin
	counter_out<= 32'h00000000;
	pwm_clk <=0;
	end	
//this always block runs on the fast 100MHz clock
always @(posedge clk) begin
	counter_out<=    counter_out + 32'h00000001;		
	if (counter_out  > 32'h00002710) begin 
		counter_out<= 32'h00000000;
		pwm_clk <= !pwm_clk;
		end
	end
	endmodule